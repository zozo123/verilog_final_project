`timescale 1ns /1ps

module add1 ( o, a, b );
  output [15:0] o;
  input [15:0] a;
  input [15:0] b;
  wire   n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163,
         n164;


  not	#(1.010) U4 ( n60, n160 );
  nor	#(1.432) U5 ( n160, n161, n162 );
  not	#(1.924) U6 ( n52, n156 );
  not	#(0.340) U7 ( n45, n152 );
  not	#(0.920) U8 ( n38, n148 );
  not	#(0.197) U9 ( n31, n144 );
  not	#(0.807) U10 ( n24, n140 );
  not	#(0.179) U11 ( n17, n136 );
  not	#(1.878) U12 ( n10, n132 );
  not	#(0.080) U13 ( n109, n107 );
  not	#(0.362) U14 ( n98, n96 );
  not	#(1.482) U15 ( n87, n85 );
  not	#(1.316) U16 ( n73, n71 );
  not	#(1.956) U17 ( n120, n118 );
  nor	#(1.449) U18 ( o[2], n50, n51 );
  and	#(0.225) U19 ( n51, n52, n53 );
  nor	#(0.646) U20 ( n50, n52, n53 );
  nand	#(0.592) U21 ( n53, n54, n55 );
  nor	#(1.762) U22 ( o[3], n43, n44 );
  and	#(0.331) U23 ( n44, n45, n46 );
  nor	#(0.068) U24 ( n43, n45, n46 );
  nand	#(0.466) U25 ( n46, n47, n48 );
  nor	#(1.628) U26 ( o[4], n36, n37 );
  and	#(0.535) U27 ( n37, n38, n39 );
  nor	#(1.244) U28 ( n36, n38, n39 );
  nand	#(1.998) U29 ( n39, n40, n41 );
  nor	#(0.570) U30 ( o[5], n29, n30 );
  and	#(0.929) U31 ( n30, n31, n32 );
  nor	#(0.902) U32 ( n29, n31, n32 );
  nand	#(0.994) U33 ( n32, n33, n34 );
  nor	#(0.210) U34 ( o[6], n22, n23 );
  and	#(0.520) U35 ( n23, n24, n25 );
  nor	#(1.417) U36 ( n22, n24, n25 );
  nand	#(1.138) U37 ( n25, n26, n27 );
  nor	#(0.057) U38 ( o[7], n15, n16 );
  and	#(0.097) U39 ( n16, n17, n18 );
  nor	#(1.457) U40 ( n15, n17, n18 );
  nand	#(0.321) U41 ( n18, n19, n20 );
  nor	#(1.763) U42 ( o[8], n8, n9 );
  and	#(1.733) U43 ( n9, n10, n11 );
  nor	#(0.729) U44 ( n8, n10, n11 );
  nand	#(0.637) U45 ( n11, n12, n13 );
  nor	#(0.388) U46 ( o[9], n1, n2 );
  and	#(1.224) U47 ( n2, n3, n4 );
  nor	#(1.914) U48 ( n1, n3, n4 );
  nand	#(0.847) U49 ( n4, n5, n6 );
  nor	#(0.253) U50 ( o[10], n121, n122 );
  and	#(0.785) U51 ( n122, n120, n123 );
  nor	#(1.825) U52 ( n121, n120, n123 );
  nand	#(1.132) U53 ( n123, n124, n125 );
  nor	#(1.940) U54 ( o[11], n110, n111 );
  and	#(0.309) U55 ( n111, n109, n112 );
  nor	#(0.882) U56 ( n110, n109, n112 );
  nand	#(0.940) U57 ( n112, n113, n114 );
  nor	#(1.989) U58 ( o[12], n99, n100 );
  and	#(0.508) U59 ( n100, n98, n101 );
  nor	#(0.936) U60 ( n99, n98, n101 );
  nand	#(1.748) U61 ( n101, n102, n103 );
  nor	#(1.877) U62 ( o[13], n88, n89 );
  and	#(0.245) U63 ( n89, n87, n90 );
  nor	#(0.530) U64 ( n88, n87, n90 );
  nand	#(1.540) U65 ( n90, n91, n92 );
  nor	#(1.818) U66 ( o[14], n77, n78 );
  and	#(1.369) U67 ( n78, n73, n79 );
  nor	#(1.639) U68 ( n77, n73, n79 );
  nand	#(0.826) U69 ( n79, n80, n81 );
  nor	#(1.965) U70 ( o[15], n64, n65 );
  and	#(1.363) U71 ( n65, n66, n67 );
  nor	#(0.969) U72 ( n64, n67, n66 );
  nand	#(1.007) U73 ( n66, n68, n69 );
  nand	#(0.569) U74 ( o[1], n57, n58 );
  or	#(1.132) U75 ( n58, n59, n60 );
  nand	#(1.863) U76 ( n57, n59, n60 );
  nand	#(0.898) U77 ( n59, n61, n62 );
  nand	#(1.649) U78 ( n3, n129, n130 );
  nand	#(0.218) U79 ( n129, a[8], n10 );
  nand	#(1.887) U80 ( n130, b[8], n131 );
  nand	#(0.226) U81 ( n131, n132, n14 );
  and	#(1.754) U82 ( n156, n157, n158 );
  nand	#(0.778) U83 ( n158, b[1], n159 );
  nand	#(0.149) U84 ( n157, a[1], n160 );
  nand	#(1.914) U85 ( n159, n63, n60 );
  and	#(0.365) U86 ( n152, n153, n154 );
  nand	#(0.627) U87 ( n153, a[2], n52 );
  nand	#(1.427) U88 ( n154, b[2], n155 );
  nand	#(1.957) U89 ( n155, n156, n56 );
  and	#(1.505) U90 ( n148, n149, n150 );
  nand	#(0.661) U91 ( n149, a[3], n45 );
  nand	#(1.154) U92 ( n150, b[3], n151 );
  nand	#(0.719) U93 ( n151, n152, n49 );
  and	#(1.118) U94 ( n144, n145, n146 );
  nand	#(0.964) U95 ( n145, a[4], n38 );
  nand	#(0.328) U96 ( n146, b[4], n147 );
  nand	#(0.438) U97 ( n147, n148, n42 );
  and	#(1.777) U98 ( n107, n115, n116 );
  nand	#(0.930) U99 ( n115, a[10], n120 );
  nand	#(0.414) U100 ( n116, b[10], n117 );
  nand	#(0.780) U101 ( n117, n118, n119 );
  and	#(1.296) U102 ( n140, n141, n142 );
  nand	#(1.692) U103 ( n141, a[5], n31 );
  nand	#(1.297) U104 ( n142, b[5], n143 );
  nand	#(1.233) U105 ( n143, n144, n35 );
  and	#(0.788) U106 ( n96, n104, n105 );
  nand	#(0.187) U107 ( n104, a[11], n109 );
  nand	#(0.346) U108 ( n105, b[11], n106 );
  nand	#(0.162) U109 ( n106, n107, n108 );
  and	#(0.747) U110 ( n136, n137, n138 );
  nand	#(1.156) U111 ( n137, a[6], n24 );
  nand	#(1.653) U112 ( n138, b[6], n139 );
  nand	#(1.338) U113 ( n139, n140, n28 );
  and	#(0.716) U114 ( n85, n93, n94 );
  nand	#(0.404) U115 ( n93, a[12], n98 );
  nand	#(1.512) U116 ( n94, b[12], n95 );
  nand	#(1.752) U117 ( n95, n96, n97 );
  and	#(1.092) U118 ( n132, n133, n134 );
  nand	#(1.621) U119 ( n133, a[7], n17 );
  nand	#(1.201) U120 ( n134, b[7], n135 );
  nand	#(1.529) U121 ( n135, n136, n21 );
  and	#(0.646) U122 ( n71, n82, n83 );
  nand	#(0.086) U123 ( n82, a[13], n87 );
  nand	#(1.122) U124 ( n83, b[13], n84 );
  nand	#(1.742) U125 ( n84, n85, n86 );
  and	#(0.302) U126 ( n118, n126, n127 );
  nand	#(1.561) U127 ( n127, b[9], n128 );
  nand	#(1.370) U128 ( n126, a[9], n3 );
  or	#(0.965) U129 ( n128, n3, a[9] );
  nand	#(0.762) U130 ( n67, n74, n75 );
  or	#(1.687) U131 ( n74, n76, b[15] );
  nand	#(0.793) U132 ( n75, b[15], n76 );
  not	#(0.348) U133 ( n76, a[15] );
  nand	#(0.512) U134 ( n55, b[2], n56 );
  nand	#(0.200) U135 ( n48, b[3], n49 );
  nand	#(1.594) U136 ( n41, b[4], n42 );
  nand	#(0.042) U137 ( n34, b[5], n35 );
  nand	#(1.795) U138 ( n27, b[6], n28 );
  nand	#(1.271) U139 ( n20, b[7], n21 );
  nand	#(1.558) U140 ( n13, b[8], n14 );
  nand	#(0.791) U141 ( n125, b[10], n119 );
  nand	#(1.097) U142 ( n114, b[11], n108 );
  nand	#(0.296) U143 ( n103, b[12], n97 );
  nand	#(0.944) U144 ( n92, b[13], n86 );
  nand	#(1.490) U145 ( n81, b[14], n72 );
  nand	#(1.719) U146 ( n62, b[1], n63 );
  nand	#(0.428) U147 ( n69, b[14], n70 );
  nand	#(0.123) U148 ( n70, n71, n72 );
  nand	#(0.525) U149 ( n68, a[14], n73 );
  not	#(0.990) U150 ( n56, a[2] );
  not	#(1.187) U151 ( n49, a[3] );
  not	#(1.012) U152 ( n42, a[4] );
  not	#(1.726) U153 ( n35, a[5] );
  not	#(1.692) U154 ( n28, a[6] );
  not	#(0.438) U155 ( n21, a[7] );
  not	#(0.375) U156 ( n14, a[8] );
  not	#(0.709) U157 ( n119, a[10] );
  not	#(0.250) U158 ( n108, a[11] );
  not	#(0.074) U159 ( n97, a[12] );
  not	#(0.045) U160 ( n86, a[13] );
  not	#(0.459) U161 ( n72, a[14] );
  nand	#(1.255) U162 ( n6, b[9], n7 );
  not	#(0.685) U163 ( n63, a[1] );
  not	#(0.140) U164 ( n161, b[0] );
  not	#(1.936) U165 ( n162, a[0] );
  nand	#(0.886) U166 ( o[0], n163, n164 );
  nand	#(1.564) U167 ( n163, a[0], n161 );
  nand	#(0.325) U168 ( n164, b[0], n162 );
  or	#(0.537) U169 ( n61, n63, b[1] );
  or	#(0.779) U170 ( n54, n56, b[2] );
  or	#(1.321) U171 ( n47, n49, b[3] );
  or	#(1.190) U172 ( n40, n42, b[4] );
  or	#(0.210) U173 ( n33, n35, b[5] );
  or	#(0.926) U174 ( n26, n28, b[6] );
  or	#(1.456) U175 ( n19, n21, b[7] );
  or	#(0.803) U176 ( n12, n14, b[8] );
  or	#(0.051) U177 ( n5, n7, b[9] );
  or	#(1.153) U178 ( n124, n119, b[10] );
  or	#(0.177) U179 ( n113, n108, b[11] );
  or	#(0.501) U180 ( n102, n97, b[12] );
  or	#(1.172) U181 ( n91, n86, b[13] );
  or	#(1.737) U182 ( n80, n72, b[14] );
  not	#(0.784) U183 ( n7, a[9] );
endmodule
