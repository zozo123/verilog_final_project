// DATA derived from module add1 !!!!!!!!!!!!!!!!
// table may be used turbosim to hold the net connectivity
// table width is 92 bits, 5x16+4+4+4
// where 5 = 1 driver + 4 loads
// where 16 = 12 + 4, 12 = cell index + bit 11 set if exist
// where 4  = pin index of driving/load cell
// next is 4 bits reflects the number of loads on net
// next is 4 bits for the current output value, set to x, R/W field
// next is 4 bits control that can be used for whatever, also R/W field
// ATTENTION : initial value of input nets/ports currently set to X !!!
000_0_84a_1_848_1_000_0_000_0_2_2_0 //    0 a[0]    |  no dpin    ,U167  pin1 ,U165  pin1 ,no load    ,no load    ,n loads 2, val x, ctl
000_0_83f_1_8b3_1_000_0_000_0_2_2_0 //    1 a[10]   |  no dpin    ,U157  pin1 ,U99   pin1 ,no load    ,no load    ,n loads 2, val x, ctl
000_0_808_1_840_1_000_0_000_0_2_2_0 //    2 a[11]   |  no dpin    ,U107  pin1 ,U158  pin1 ,no load    ,no load    ,n loads 2, val x, ctl
000_0_811_1_841_1_000_0_000_0_2_2_0 //    3 a[12]   |  no dpin    ,U115  pin1 ,U159  pin1 ,no load    ,no load    ,n loads 2, val x, ctl
000_0_843_1_81a_1_000_0_000_0_2_2_0 //    4 a[13]   |  no dpin    ,U160  pin1 ,U123  pin1 ,no load    ,no load    ,n loads 2, val x, ctl
000_0_836_1_844_1_000_0_000_0_2_2_0 //    5 a[14]   |  no dpin    ,U149  pin1 ,U161  pin1 ,no load    ,no load    ,n loads 2, val x, ctl
000_0_825_1_000_0_000_0_000_0_1_2_0 //    6 a[15]   |  no dpin    ,U133  pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
000_0_846_1_8a3_1_000_0_000_0_2_2_0 //    7 a[1]    |  no dpin    ,U163  pin1 ,U84   pin1 ,no load    ,no load    ,n loads 2, val x, ctl
000_0_8a6_1_838_1_000_0_000_0_2_2_0 //    8 a[2]    |  no dpin    ,U87   pin1 ,U150  pin1 ,no load    ,no load    ,n loads 2, val x, ctl
000_0_839_1_8ab_1_000_0_000_0_2_2_0 //    9 a[3]    |  no dpin    ,U151  pin1 ,U91   pin1 ,no load    ,no load    ,n loads 2, val x, ctl
000_0_83a_1_8af_1_000_0_000_0_2_2_0 //   10 a[4]    |  no dpin    ,U152  pin1 ,U95   pin1 ,no load    ,no load    ,n loads 2, val x, ctl
000_0_83b_1_804_1_000_0_000_0_2_2_0 //   11 a[5]    |  no dpin    ,U153  pin1 ,U103  pin1 ,no load    ,no load    ,n loads 2, val x, ctl
000_0_83c_1_80d_1_000_0_000_0_2_2_0 //   12 a[6]    |  no dpin    ,U154  pin1 ,U111  pin1 ,no load    ,no load    ,n loads 2, val x, ctl
000_0_815_1_83d_1_000_0_000_0_2_2_0 //   13 a[7]    |  no dpin    ,U119  pin1 ,U155  pin1 ,no load    ,no load    ,n loads 2, val x, ctl
000_0_83e_1_89d_1_000_0_000_0_2_2_0 //   14 a[8]    |  no dpin    ,U156  pin1 ,U79   pin1 ,no load    ,no load    ,n loads 2, val x, ctl
000_0_820_2_85c_1_81f_1_000_0_3_2_0 //   15 a[9]    |  no dpin    ,U129  pin2 ,U183  pin1 ,U128  pin1 ,no load    ,n loads 3, val x, ctl
000_0_847_1_84b_1_000_0_000_0_2_2_0 //   16 b[0]    |  no dpin    ,U164  pin1 ,U168  pin1 ,no load    ,no load    ,n loads 2, val x, ctl
000_0_856_2_82e_1_801_1_000_0_3_2_0 //   17 b[10]   |  no dpin    ,U178  pin2 ,U141  pin1 ,U100  pin1 ,no load    ,n loads 3, val x, ctl
000_0_857_2_809_1_82f_1_000_0_3_2_0 //   18 b[11]   |  no dpin    ,U179  pin2 ,U108  pin1 ,U142  pin1 ,no load    ,n loads 3, val x, ctl
000_0_830_1_812_1_859_2_000_0_3_2_0 //   19 b[12]   |  no dpin    ,U143  pin1 ,U116  pin1 ,U180  pin2 ,no load    ,n loads 3, val x, ctl
000_0_81b_1_85a_2_831_1_000_0_3_2_0 //   20 b[13]   |  no dpin    ,U124  pin1 ,U181  pin2 ,U144  pin1 ,no load    ,n loads 3, val x, ctl
000_0_85b_2_834_1_832_1_000_0_3_2_0 //   21 b[14]   |  no dpin    ,U182  pin2 ,U147  pin1 ,U145  pin1 ,no load    ,n loads 3, val x, ctl
000_0_823_2_824_1_000_0_000_0_2_2_0 //   22 b[15]   |  no dpin    ,U131  pin2 ,U132  pin1 ,no load    ,no load    ,n loads 2, val x, ctl
000_0_833_1_84c_2_8a2_1_000_0_3_2_0 //   23 b[1]    |  no dpin    ,U146  pin1 ,U169  pin2 ,U83   pin1 ,no load    ,n loads 3, val x, ctl
000_0_8a7_1_84e_2_826_1_000_0_3_2_0 //   24 b[2]    |  no dpin    ,U88   pin1 ,U170  pin2 ,U134  pin1 ,no load    ,n loads 3, val x, ctl
000_0_827_1_84f_2_8ac_1_000_0_3_2_0 //   25 b[3]    |  no dpin    ,U135  pin1 ,U171  pin2 ,U92   pin1 ,no load    ,n loads 3, val x, ctl
000_0_850_2_828_1_8b0_1_000_0_3_2_0 //   26 b[4]    |  no dpin    ,U172  pin2 ,U136  pin1 ,U96   pin1 ,no load    ,n loads 3, val x, ctl
000_0_805_1_851_2_829_1_000_0_3_2_0 //   27 b[5]    |  no dpin    ,U104  pin1 ,U173  pin2 ,U137  pin1 ,no load    ,n loads 3, val x, ctl
000_0_82a_1_852_2_80e_1_000_0_3_2_0 //   28 b[6]    |  no dpin    ,U138  pin1 ,U174  pin2 ,U112  pin1 ,no load    ,n loads 3, val x, ctl
000_0_82b_1_853_2_817_1_000_0_3_2_0 //   29 b[7]    |  no dpin    ,U139  pin1 ,U175  pin2 ,U120  pin1 ,no load    ,n loads 3, val x, ctl
000_0_854_2_89f_1_82d_1_000_0_3_2_0 //   30 b[8]    |  no dpin    ,U176  pin2 ,U80   pin1 ,U140  pin1 ,no load    ,n loads 3, val x, ctl
000_0_845_1_81e_1_855_2_000_0_3_2_0 //   31 b[9]    |  no dpin    ,U162  pin1 ,U127  pin1 ,U177  pin2 ,no load    ,n loads 3, val x, ctl
87b_0_879_1_000_0_000_0_000_0_1_2_0 //   32 n1      |  U48   pin0 ,U46   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
816_0_877_1_89d_2_876_1_000_0_3_2_0 //   33 n10     |  U12   pin0 ,U44   pin1 ,U79   pin2 ,U43   pin1 ,no load    ,n loads 3, val x, ctl
887_0_886_2_000_0_000_0_000_0_1_2_0 //   34 n100    |  U59   pin0 ,U58   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
88a_0_887_2_889_2_000_0_000_0_2_2_0 //   35 n101    |  U61   pin0 ,U59   pin2 ,U60   pin2 ,no load    ,no load    ,n loads 2, val x, ctl
859_0_88a_1_000_0_000_0_000_0_1_2_0 //   36 n102    |  U180  pin0 ,U61   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
830_0_88a_2_000_0_000_0_000_0_1_2_0 //   37 n103    |  U143  pin0 ,U61   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
808_0_807_1_000_0_000_0_000_0_1_2_0 //   38 n104    |  U107  pin0 ,U106  pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
809_0_807_2_000_0_000_0_000_0_1_2_0 //   39 n105    |  U108  pin0 ,U106  pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
80a_0_809_2_000_0_000_0_000_0_1_2_0 //   40 n106    |  U109  pin0 ,U108  pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
8b2_0_80a_1_821_1_000_0_000_0_2_2_0 //   41 n107    |  U98   pin0 ,U109  pin1 ,U13   pin1 ,no load    ,no load    ,n loads 2, val x, ctl
840_0_82f_2_80a_2_857_1_000_0_3_2_0 //   42 n108    |  U158  pin0 ,U142  pin2 ,U109  pin2 ,U179  pin1 ,no load    ,n loads 3, val x, ctl
821_0_884_1_883_1_808_2_000_0_3_2_0 //   43 n109    |  U13   pin0 ,U56   pin1 ,U55   pin1 ,U107  pin2 ,no load    ,n loads 3, val x, ctl
878_0_876_2_877_2_000_0_000_0_2_2_0 //   44 n11     |  U45   pin0 ,U43   pin2 ,U44   pin2 ,no load    ,no load    ,n loads 2, val x, ctl
884_0_882_1_000_0_000_0_000_0_1_2_0 //   45 n110    |  U56   pin0 ,U54   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
883_0_882_2_000_0_000_0_000_0_1_2_0 //   46 n111    |  U55   pin0 ,U54   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
885_0_884_2_883_2_000_0_000_0_2_2_0 //   47 n112    |  U57   pin0 ,U56   pin2 ,U55   pin2 ,no load    ,no load    ,n loads 2, val x, ctl
857_0_885_1_000_0_000_0_000_0_1_2_0 //   48 n113    |  U179  pin0 ,U57   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
82f_0_885_2_000_0_000_0_000_0_1_2_0 //   49 n114    |  U142  pin0 ,U57   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
8b3_0_8b2_1_000_0_000_0_000_0_1_2_0 //   50 n115    |  U99   pin0 ,U98   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
801_0_8b2_2_000_0_000_0_000_0_1_2_0 //   51 n116    |  U100  pin0 ,U98   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
802_0_801_2_000_0_000_0_000_0_1_2_0 //   52 n117    |  U101  pin0 ,U100  pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
81d_0_802_1_84d_1_000_0_000_0_2_2_0 //   53 n118    |  U126  pin0 ,U101  pin1 ,U17   pin1 ,no load    ,no load    ,n loads 2, val x, ctl
83f_0_82e_2_856_1_802_2_000_0_3_2_0 //   54 n119    |  U157  pin0 ,U141  pin2 ,U178  pin1 ,U101  pin2 ,no load    ,n loads 3, val x, ctl
854_0_878_1_000_0_000_0_000_0_1_2_0 //   55 n12     |  U176  pin0 ,U45   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
84d_0_8b3_2_880_1_87f_1_000_0_3_2_0 //   56 n120    |  U17   pin0 ,U99   pin2 ,U52   pin1 ,U51   pin1 ,no load    ,n loads 3, val x, ctl
880_0_87e_1_000_0_000_0_000_0_1_2_0 //   57 n121    |  U52   pin0 ,U50   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
87f_0_87e_2_000_0_000_0_000_0_1_2_0 //   58 n122    |  U51   pin0 ,U50   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
881_0_880_2_87f_2_000_0_000_0_2_2_0 //   59 n123    |  U53   pin0 ,U52   pin2 ,U51   pin2 ,no load    ,no load    ,n loads 2, val x, ctl
856_0_881_1_000_0_000_0_000_0_1_2_0 //   60 n124    |  U178  pin0 ,U53   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
82e_0_881_2_000_0_000_0_000_0_1_2_0 //   61 n125    |  U141  pin0 ,U53   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
81f_0_81d_1_000_0_000_0_000_0_1_2_0 //   62 n126    |  U128  pin0 ,U126  pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
81e_0_81d_2_000_0_000_0_000_0_1_2_0 //   63 n127    |  U127  pin0 ,U126  pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
820_0_81e_2_000_0_000_0_000_0_1_2_0 //   64 n128    |  U129  pin0 ,U127  pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
89d_0_89c_1_000_0_000_0_000_0_1_2_0 //   65 n129    |  U79   pin0 ,U78   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
82d_0_878_2_000_0_000_0_000_0_1_2_0 //   66 n13     |  U140  pin0 ,U45   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
89f_0_89c_2_000_0_000_0_000_0_1_2_0 //   67 n130    |  U80   pin0 ,U78   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
8a0_0_89f_2_000_0_000_0_000_0_1_2_0 //   68 n131    |  U81   pin0 ,U80   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
814_0_816_1_8a0_1_000_0_000_0_2_2_0 //   69 n132    |  U118  pin0 ,U12   pin1 ,U81   pin1 ,no load    ,no load    ,n loads 2, val x, ctl
815_0_814_1_000_0_000_0_000_0_1_2_0 //   70 n133    |  U119  pin0 ,U118  pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
817_0_814_2_000_0_000_0_000_0_1_2_0 //   71 n134    |  U120  pin0 ,U118  pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
818_0_817_2_000_0_000_0_000_0_1_2_0 //   72 n135    |  U121  pin0 ,U120  pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
80c_0_818_1_80b_1_000_0_000_0_2_2_0 //   73 n136    |  U110  pin0 ,U121  pin1 ,U11   pin1 ,no load    ,no load    ,n loads 2, val x, ctl
80d_0_80c_1_000_0_000_0_000_0_1_2_0 //   74 n137    |  U111  pin0 ,U110  pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
80e_0_80c_2_000_0_000_0_000_0_1_2_0 //   75 n138    |  U112  pin0 ,U110  pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
80f_0_80e_2_000_0_000_0_000_0_1_2_0 //   76 n139    |  U113  pin0 ,U112  pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
83e_0_8a0_2_854_1_82d_2_000_0_3_2_0 //   77 n14     |  U156  pin0 ,U81   pin2 ,U176  pin1 ,U140  pin2 ,no load    ,n loads 3, val x, ctl
803_0_80f_1_800_1_000_0_000_0_2_2_0 //   78 n140    |  U102  pin0 ,U113  pin1 ,U10   pin1 ,no load    ,no load    ,n loads 2, val x, ctl
804_0_803_1_000_0_000_0_000_0_1_2_0 //   79 n141    |  U103  pin0 ,U102  pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
805_0_803_2_000_0_000_0_000_0_1_2_0 //   80 n142    |  U104  pin0 ,U102  pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
806_0_805_2_000_0_000_0_000_0_1_2_0 //   81 n143    |  U105  pin0 ,U104  pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
8ae_0_806_1_8a9_1_000_0_000_0_2_2_0 //   82 n144    |  U94   pin0 ,U105  pin1 ,U9    pin1 ,no load    ,no load    ,n loads 2, val x, ctl
8af_0_8ae_1_000_0_000_0_000_0_1_2_0 //   83 n145    |  U95   pin0 ,U94   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
8b0_0_8ae_2_000_0_000_0_000_0_1_2_0 //   84 n146    |  U96   pin0 ,U94   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
8b1_0_8b0_2_000_0_000_0_000_0_1_2_0 //   85 n147    |  U97   pin0 ,U96   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
8aa_0_8b1_1_89e_1_000_0_000_0_2_2_0 //   86 n148    |  U90   pin0 ,U97   pin1 ,U8    pin1 ,no load    ,no load    ,n loads 2, val x, ctl
8ab_0_8aa_1_000_0_000_0_000_0_1_2_0 //   87 n149    |  U91   pin0 ,U90   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
873_0_870_1_000_0_000_0_000_0_1_2_0 //   88 n15     |  U40   pin0 ,U38   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
8ac_0_8aa_2_000_0_000_0_000_0_1_2_0 //   89 n150    |  U92   pin0 ,U90   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
8ad_0_8ac_2_000_0_000_0_000_0_1_2_0 //   90 n151    |  U93   pin0 ,U92   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
8a5_0_893_1_8ad_1_000_0_000_0_2_2_0 //   91 n152    |  U86   pin0 ,U7    pin1 ,U93   pin1 ,no load    ,no load    ,n loads 2, val x, ctl
8a6_0_8a5_1_000_0_000_0_000_0_1_2_0 //   92 n153    |  U87   pin0 ,U86   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
8a7_0_8a5_2_000_0_000_0_000_0_1_2_0 //   93 n154    |  U88   pin0 ,U86   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
8a8_0_8a7_2_000_0_000_0_000_0_1_2_0 //   94 n155    |  U89   pin0 ,U88   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
8a1_0_888_1_8a8_1_000_0_000_0_2_2_0 //   95 n156    |  U82   pin0 ,U6    pin1 ,U89   pin1 ,no load    ,no load    ,n loads 2, val x, ctl
8a3_0_8a1_1_000_0_000_0_000_0_1_2_0 //   96 n157    |  U84   pin0 ,U82   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
8a2_0_8a1_2_000_0_000_0_000_0_1_2_0 //   97 n158    |  U83   pin0 ,U82   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
8a4_0_8a2_2_000_0_000_0_000_0_1_2_0 //   98 n159    |  U85   pin0 ,U83   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
871_0_870_2_000_0_000_0_000_0_1_2_0 //   99 n16     |  U39   pin0 ,U38   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
87d_0_872_1_8a3_2_000_0_000_0_2_2_0 //  100 n160    |  U5    pin0 ,U4    pin1 ,U84   pin2 ,no load    ,no load    ,n loads 2, val x, ctl
847_0_84a_2_87d_1_000_0_000_0_2_2_0 //  101 n161    |  U164  pin0 ,U167  pin2 ,U5    pin1 ,no load    ,no load    ,n loads 2, val x, ctl
848_0_87d_2_84b_2_000_0_000_0_2_2_0 //  102 n162    |  U165  pin0 ,U5    pin2 ,U168  pin2 ,no load    ,no load    ,n loads 2, val x, ctl
84a_0_849_1_000_0_000_0_000_0_1_2_0 //  103 n163    |  U167  pin0 ,U166  pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
84b_0_849_2_000_0_000_0_000_0_1_2_0 //  104 n164    |  U168  pin0 ,U166  pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
80b_0_871_1_873_1_815_2_000_0_3_2_0 //  105 n17     |  U11   pin0 ,U39   pin1 ,U40   pin1 ,U119  pin2 ,no load    ,n loads 3, val x, ctl
874_0_873_2_871_2_000_0_000_0_2_2_0 //  106 n18     |  U41   pin0 ,U40   pin2 ,U39   pin2 ,no load    ,no load    ,n loads 2, val x, ctl
853_0_874_1_000_0_000_0_000_0_1_2_0 //  107 n19     |  U175  pin0 ,U41   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
87a_0_879_2_000_0_000_0_000_0_1_2_0 //  108 n2      |  U47   pin0 ,U46   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
82b_0_874_2_000_0_000_0_000_0_1_2_0 //  109 n20     |  U139  pin0 ,U41   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
83d_0_82b_2_853_1_818_2_000_0_3_2_0 //  110 n21     |  U155  pin0 ,U139  pin2 ,U175  pin1 ,U121  pin2 ,no load    ,n loads 3, val x, ctl
86e_0_86c_1_000_0_000_0_000_0_1_2_0 //  111 n22     |  U36   pin0 ,U34   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
86d_0_86c_2_000_0_000_0_000_0_1_2_0 //  112 n23     |  U35   pin0 ,U34   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
800_0_80d_2_86e_1_86d_1_000_0_3_2_0 //  113 n24     |  U10   pin0 ,U111  pin2 ,U36   pin1 ,U35   pin1 ,no load    ,n loads 3, val x, ctl
86f_0_86e_2_86d_2_000_0_000_0_2_2_0 //  114 n25     |  U37   pin0 ,U36   pin2 ,U35   pin2 ,no load    ,no load    ,n loads 2, val x, ctl
852_0_86f_1_000_0_000_0_000_0_1_2_0 //  115 n26     |  U174  pin0 ,U37   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
82a_0_86f_2_000_0_000_0_000_0_1_2_0 //  116 n27     |  U138  pin0 ,U37   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
83c_0_852_1_80f_2_82a_2_000_0_3_2_0 //  117 n28     |  U154  pin0 ,U174  pin1 ,U113  pin2 ,U138  pin2 ,no load    ,n loads 3, val x, ctl
86a_0_868_1_000_0_000_0_000_0_1_2_0 //  118 n29     |  U32   pin0 ,U30   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
89c_0_820_1_87b_1_87a_1_81f_2_4_2_0 //  119 n3      |  U78   pin0 ,U129  pin1 ,U48   pin1 ,U47   pin1 ,U128  pin2 ,n loads 4, val x, ctl
869_0_868_2_000_0_000_0_000_0_1_2_0 //  120 n30     |  U31   pin0 ,U30   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
8a9_0_86a_1_869_1_804_2_000_0_3_2_0 //  121 n31     |  U9    pin0 ,U32   pin1 ,U31   pin1 ,U103  pin2 ,no load    ,n loads 3, val x, ctl
86b_0_869_2_86a_2_000_0_000_0_2_2_0 //  122 n32     |  U33   pin0 ,U31   pin2 ,U32   pin2 ,no load    ,no load    ,n loads 2, val x, ctl
851_0_86b_1_000_0_000_0_000_0_1_2_0 //  123 n33     |  U173  pin0 ,U33   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
829_0_86b_2_000_0_000_0_000_0_1_2_0 //  124 n34     |  U137  pin0 ,U33   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
83b_0_851_1_829_2_806_2_000_0_3_2_0 //  125 n35     |  U153  pin0 ,U173  pin1 ,U137  pin2 ,U105  pin2 ,no load    ,n loads 3, val x, ctl
866_0_864_1_000_0_000_0_000_0_1_2_0 //  126 n36     |  U28   pin0 ,U26   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
865_0_864_2_000_0_000_0_000_0_1_2_0 //  127 n37     |  U27   pin0 ,U26   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
89e_0_865_1_8af_2_866_1_000_0_3_2_0 //  128 n38     |  U8    pin0 ,U27   pin1 ,U95   pin2 ,U28   pin1 ,no load    ,n loads 3, val x, ctl
867_0_866_2_865_2_000_0_000_0_2_2_0 //  129 n39     |  U29   pin0 ,U28   pin2 ,U27   pin2 ,no load    ,no load    ,n loads 2, val x, ctl
87c_0_87a_2_87b_2_000_0_000_0_2_2_0 //  130 n4      |  U49   pin0 ,U47   pin2 ,U48   pin2 ,no load    ,no load    ,n loads 2, val x, ctl
850_0_867_1_000_0_000_0_000_0_1_2_0 //  131 n40     |  U172  pin0 ,U29   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
828_0_867_2_000_0_000_0_000_0_1_2_0 //  132 n41     |  U136  pin0 ,U29   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
83a_0_850_1_8b1_2_828_2_000_0_3_2_0 //  133 n42     |  U152  pin0 ,U172  pin1 ,U97   pin2 ,U136  pin2 ,no load    ,n loads 3, val x, ctl
862_0_860_1_000_0_000_0_000_0_1_2_0 //  134 n43     |  U24   pin0 ,U22   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
861_0_860_2_000_0_000_0_000_0_1_2_0 //  135 n44     |  U23   pin0 ,U22   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
893_0_862_1_8ab_2_861_1_000_0_3_2_0 //  136 n45     |  U7    pin0 ,U24   pin1 ,U91   pin2 ,U23   pin1 ,no load    ,n loads 3, val x, ctl
863_0_862_2_861_2_000_0_000_0_2_2_0 //  137 n46     |  U25   pin0 ,U24   pin2 ,U23   pin2 ,no load    ,no load    ,n loads 2, val x, ctl
84f_0_863_1_000_0_000_0_000_0_1_2_0 //  138 n47     |  U171  pin0 ,U25   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
827_0_863_2_000_0_000_0_000_0_1_2_0 //  139 n48     |  U135  pin0 ,U25   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
839_0_8ad_2_827_2_84f_1_000_0_3_2_0 //  140 n49     |  U151  pin0 ,U93   pin2 ,U135  pin2 ,U171  pin1 ,no load    ,n loads 3, val x, ctl
855_0_87c_1_000_0_000_0_000_0_1_2_0 //  141 n5      |  U177  pin0 ,U49   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
85e_0_858_1_000_0_000_0_000_0_1_2_0 //  142 n50     |  U20   pin0 ,U18   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
85d_0_858_2_000_0_000_0_000_0_1_2_0 //  143 n51     |  U19   pin0 ,U18   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
888_0_85d_1_85e_1_8a6_2_000_0_3_2_0 //  144 n52     |  U6    pin0 ,U19   pin1 ,U20   pin1 ,U87   pin2 ,no load    ,n loads 3, val x, ctl
85f_0_85e_2_85d_2_000_0_000_0_2_2_0 //  145 n53     |  U21   pin0 ,U20   pin2 ,U19   pin2 ,no load    ,no load    ,n loads 2, val x, ctl
84e_0_85f_1_000_0_000_0_000_0_1_2_0 //  146 n54     |  U170  pin0 ,U21   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
826_0_85f_2_000_0_000_0_000_0_1_2_0 //  147 n55     |  U134  pin0 ,U21   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
838_0_84e_1_826_2_8a8_2_000_0_3_2_0 //  148 n56     |  U150  pin0 ,U170  pin1 ,U134  pin2 ,U89   pin2 ,no load    ,n loads 3, val x, ctl
89a_0_898_1_000_0_000_0_000_0_1_2_0 //  149 n57     |  U76   pin0 ,U74   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
899_0_898_2_000_0_000_0_000_0_1_2_0 //  150 n58     |  U75   pin0 ,U74   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
89b_0_89a_1_899_1_000_0_000_0_2_2_0 //  151 n59     |  U77   pin0 ,U76   pin1 ,U75   pin1 ,no load    ,no load    ,n loads 2, val x, ctl
845_0_87c_2_000_0_000_0_000_0_1_2_0 //  152 n6      |  U162  pin0 ,U49   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
872_0_899_2_8a4_2_89a_2_000_0_3_2_0 //  153 n60     |  U4    pin0 ,U75   pin2 ,U85   pin2 ,U76   pin2 ,no load    ,n loads 3, val x, ctl
84c_0_89b_1_000_0_000_0_000_0_1_2_0 //  154 n61     |  U169  pin0 ,U77   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
833_0_89b_2_000_0_000_0_000_0_1_2_0 //  155 n62     |  U146  pin0 ,U77   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
846_0_8a4_1_84c_1_833_2_000_0_3_2_0 //  156 n63     |  U163  pin0 ,U85   pin1 ,U169  pin1 ,U146  pin2 ,no load    ,n loads 3, val x, ctl
896_0_894_1_000_0_000_0_000_0_1_2_0 //  157 n64     |  U72   pin0 ,U70   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
895_0_894_2_000_0_000_0_000_0_1_2_0 //  158 n65     |  U71   pin0 ,U70   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
897_0_895_1_896_2_000_0_000_0_2_2_0 //  159 n66     |  U73   pin0 ,U71   pin1 ,U72   pin2 ,no load    ,no load    ,n loads 2, val x, ctl
822_0_896_1_895_2_000_0_000_0_2_2_0 //  160 n67     |  U130  pin0 ,U72   pin1 ,U71   pin2 ,no load    ,no load    ,n loads 2, val x, ctl
836_0_897_1_000_0_000_0_000_0_1_2_0 //  161 n68     |  U149  pin0 ,U73   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
834_0_897_2_000_0_000_0_000_0_1_2_0 //  162 n69     |  U147  pin0 ,U73   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
85c_0_855_1_845_2_000_0_000_0_2_2_0 //  163 n7      |  U183  pin0 ,U177  pin1 ,U162  pin2 ,no load    ,no load    ,n loads 2, val x, ctl
835_0_834_2_000_0_000_0_000_0_1_2_0 //  164 n70     |  U148  pin0 ,U147  pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
819_0_842_1_835_1_000_0_000_0_2_2_0 //  165 n71     |  U122  pin0 ,U16   pin1 ,U148  pin1 ,no load    ,no load    ,n loads 2, val x, ctl
844_0_85b_1_832_2_835_2_000_0_3_2_0 //  166 n72     |  U161  pin0 ,U182  pin1 ,U145  pin2 ,U148  pin2 ,no load    ,n loads 3, val x, ctl
842_0_836_2_891_1_890_1_000_0_3_2_0 //  167 n73     |  U16   pin0 ,U149  pin2 ,U68   pin1 ,U67   pin1 ,no load    ,n loads 3, val x, ctl
823_0_822_1_000_0_000_0_000_0_1_2_0 //  168 n74     |  U131  pin0 ,U130  pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
824_0_822_2_000_0_000_0_000_0_1_2_0 //  169 n75     |  U132  pin0 ,U130  pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
825_0_824_2_823_1_000_0_000_0_2_2_0 //  170 n76     |  U133  pin0 ,U132  pin2 ,U131  pin1 ,no load    ,no load    ,n loads 2, val x, ctl
891_0_88f_1_000_0_000_0_000_0_1_2_0 //  171 n77     |  U68   pin0 ,U66   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
890_0_88f_2_000_0_000_0_000_0_1_2_0 //  172 n78     |  U67   pin0 ,U66   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
892_0_890_2_891_2_000_0_000_0_2_2_0 //  173 n79     |  U69   pin0 ,U67   pin2 ,U68   pin2 ,no load    ,no load    ,n loads 2, val x, ctl
877_0_875_1_000_0_000_0_000_0_1_2_0 //  174 n8      |  U44   pin0 ,U42   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
85b_0_892_1_000_0_000_0_000_0_1_2_0 //  175 n80     |  U182  pin0 ,U69   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
832_0_892_2_000_0_000_0_000_0_1_2_0 //  176 n81     |  U145  pin0 ,U69   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
81a_0_819_1_000_0_000_0_000_0_1_2_0 //  177 n82     |  U123  pin0 ,U122  pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
81b_0_819_2_000_0_000_0_000_0_1_2_0 //  178 n83     |  U124  pin0 ,U122  pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
81c_0_81b_2_000_0_000_0_000_0_1_2_0 //  179 n84     |  U125  pin0 ,U124  pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
810_0_81c_1_837_1_000_0_000_0_2_2_0 //  180 n85     |  U114  pin0 ,U125  pin1 ,U15   pin1 ,no load    ,no load    ,n loads 2, val x, ctl
843_0_81c_2_831_2_85a_1_000_0_3_2_0 //  181 n86     |  U160  pin0 ,U125  pin2 ,U144  pin2 ,U181  pin1 ,no load    ,n loads 3, val x, ctl
837_0_81a_2_88d_1_88c_1_000_0_3_2_0 //  182 n87     |  U15   pin0 ,U123  pin2 ,U64   pin1 ,U63   pin1 ,no load    ,n loads 3, val x, ctl
88d_0_88b_1_000_0_000_0_000_0_1_2_0 //  183 n88     |  U64   pin0 ,U62   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
88c_0_88b_2_000_0_000_0_000_0_1_2_0 //  184 n89     |  U63   pin0 ,U62   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
876_0_875_2_000_0_000_0_000_0_1_2_0 //  185 n9      |  U43   pin0 ,U42   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
88e_0_88d_2_88c_2_000_0_000_0_2_2_0 //  186 n90     |  U65   pin0 ,U64   pin2 ,U63   pin2 ,no load    ,no load    ,n loads 2, val x, ctl
85a_0_88e_1_000_0_000_0_000_0_1_2_0 //  187 n91     |  U181  pin0 ,U65   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
831_0_88e_2_000_0_000_0_000_0_1_2_0 //  188 n92     |  U144  pin0 ,U65   pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
811_0_810_1_000_0_000_0_000_0_1_2_0 //  189 n93     |  U115  pin0 ,U114  pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
812_0_810_2_000_0_000_0_000_0_1_2_0 //  190 n94     |  U116  pin0 ,U114  pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
813_0_812_2_000_0_000_0_000_0_1_2_0 //  191 n95     |  U117  pin0 ,U116  pin2 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
807_0_82c_1_813_1_000_0_000_0_2_2_0 //  192 n96     |  U106  pin0 ,U14   pin1 ,U117  pin1 ,no load    ,no load    ,n loads 2, val x, ctl
841_0_830_2_859_1_813_2_000_0_3_2_0 //  193 n97     |  U159  pin0 ,U143  pin2 ,U180  pin1 ,U117  pin2 ,no load    ,n loads 3, val x, ctl
82c_0_811_2_887_1_889_1_000_0_3_2_0 //  194 n98     |  U14   pin0 ,U115  pin2 ,U59   pin1 ,U60   pin1 ,no load    ,n loads 3, val x, ctl
889_0_886_1_000_0_000_0_000_0_1_2_0 //  195 n99     |  U60   pin0 ,U58   pin1 ,no load    ,no load    ,no load    ,n loads 1, val x, ctl
849_0_000_0_000_0_000_0_000_0_0_2_0 //  196 o[0]    |  U166  pin0 ,no load    ,no load    ,no load    ,no load    ,n loads 0, val x, ctl
87e_0_000_0_000_0_000_0_000_0_0_2_0 //  197 o[10]   |  U50   pin0 ,no load    ,no load    ,no load    ,no load    ,n loads 0, val x, ctl
882_0_000_0_000_0_000_0_000_0_0_2_0 //  198 o[11]   |  U54   pin0 ,no load    ,no load    ,no load    ,no load    ,n loads 0, val x, ctl
886_0_000_0_000_0_000_0_000_0_0_2_0 //  199 o[12]   |  U58   pin0 ,no load    ,no load    ,no load    ,no load    ,n loads 0, val x, ctl
88b_0_000_0_000_0_000_0_000_0_0_2_0 //  200 o[13]   |  U62   pin0 ,no load    ,no load    ,no load    ,no load    ,n loads 0, val x, ctl
88f_0_000_0_000_0_000_0_000_0_0_2_0 //  201 o[14]   |  U66   pin0 ,no load    ,no load    ,no load    ,no load    ,n loads 0, val x, ctl
894_0_000_0_000_0_000_0_000_0_0_2_0 //  202 o[15]   |  U70   pin0 ,no load    ,no load    ,no load    ,no load    ,n loads 0, val x, ctl
898_0_000_0_000_0_000_0_000_0_0_2_0 //  203 o[1]    |  U74   pin0 ,no load    ,no load    ,no load    ,no load    ,n loads 0, val x, ctl
858_0_000_0_000_0_000_0_000_0_0_2_0 //  204 o[2]    |  U18   pin0 ,no load    ,no load    ,no load    ,no load    ,n loads 0, val x, ctl
860_0_000_0_000_0_000_0_000_0_0_2_0 //  205 o[3]    |  U22   pin0 ,no load    ,no load    ,no load    ,no load    ,n loads 0, val x, ctl
864_0_000_0_000_0_000_0_000_0_0_2_0 //  206 o[4]    |  U26   pin0 ,no load    ,no load    ,no load    ,no load    ,n loads 0, val x, ctl
868_0_000_0_000_0_000_0_000_0_0_2_0 //  207 o[5]    |  U30   pin0 ,no load    ,no load    ,no load    ,no load    ,n loads 0, val x, ctl
86c_0_000_0_000_0_000_0_000_0_0_2_0 //  208 o[6]    |  U34   pin0 ,no load    ,no load    ,no load    ,no load    ,n loads 0, val x, ctl
870_0_000_0_000_0_000_0_000_0_0_2_0 //  209 o[7]    |  U38   pin0 ,no load    ,no load    ,no load    ,no load    ,n loads 0, val x, ctl
875_0_000_0_000_0_000_0_000_0_0_2_0 //  210 o[8]    |  U42   pin0 ,no load    ,no load    ,no load    ,no load    ,n loads 0, val x, ctl
879_0_000_0_000_0_000_0_000_0_0_2_0 //  211 o[9]    |  U46   pin0 ,no load    ,no load    ,no load    ,no load    ,n loads 0, val x, ctl
