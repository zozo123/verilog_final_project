// DATA derived from module add1 !!!!!!!!!!!!!!!!
// table used by testbench to translate out_records
// from turbosim to screen prints with time, value and net name
615b305d20202020202020202020202020202020 //  net index:     0, net name:     a[0]                 input
615b31305d202020202020202020202020202020 //  net index:     1, net name:     a[10]                input
615b31315d202020202020202020202020202020 //  net index:     2, net name:     a[11]                input
615b31325d202020202020202020202020202020 //  net index:     3, net name:     a[12]                input
615b31335d202020202020202020202020202020 //  net index:     4, net name:     a[13]                input
615b31345d202020202020202020202020202020 //  net index:     5, net name:     a[14]                input
615b31355d202020202020202020202020202020 //  net index:     6, net name:     a[15]                input
615b315d20202020202020202020202020202020 //  net index:     7, net name:     a[1]                 input
615b325d20202020202020202020202020202020 //  net index:     8, net name:     a[2]                 input
615b335d20202020202020202020202020202020 //  net index:     9, net name:     a[3]                 input
615b345d20202020202020202020202020202020 //  net index:    10, net name:     a[4]                 input
615b355d20202020202020202020202020202020 //  net index:    11, net name:     a[5]                 input
615b365d20202020202020202020202020202020 //  net index:    12, net name:     a[6]                 input
615b375d20202020202020202020202020202020 //  net index:    13, net name:     a[7]                 input
615b385d20202020202020202020202020202020 //  net index:    14, net name:     a[8]                 input
615b395d20202020202020202020202020202020 //  net index:    15, net name:     a[9]                 input
625b305d20202020202020202020202020202020 //  net index:    16, net name:     b[0]                 input
625b31305d202020202020202020202020202020 //  net index:    17, net name:     b[10]                input
625b31315d202020202020202020202020202020 //  net index:    18, net name:     b[11]                input
625b31325d202020202020202020202020202020 //  net index:    19, net name:     b[12]                input
625b31335d202020202020202020202020202020 //  net index:    20, net name:     b[13]                input
625b31345d202020202020202020202020202020 //  net index:    21, net name:     b[14]                input
625b31355d202020202020202020202020202020 //  net index:    22, net name:     b[15]                input
625b315d20202020202020202020202020202020 //  net index:    23, net name:     b[1]                 input
625b325d20202020202020202020202020202020 //  net index:    24, net name:     b[2]                 input
625b335d20202020202020202020202020202020 //  net index:    25, net name:     b[3]                 input
625b345d20202020202020202020202020202020 //  net index:    26, net name:     b[4]                 input
625b355d20202020202020202020202020202020 //  net index:    27, net name:     b[5]                 input
625b365d20202020202020202020202020202020 //  net index:    28, net name:     b[6]                 input
625b375d20202020202020202020202020202020 //  net index:    29, net name:     b[7]                 input
625b385d20202020202020202020202020202020 //  net index:    30, net name:     b[8]                 input
625b395d20202020202020202020202020202020 //  net index:    31, net name:     b[9]                 input
6e31202020202020202020202020202020202020 //  net index:    32, net name:     n1                   
6e31302020202020202020202020202020202020 //  net index:    33, net name:     n10                  
6e31303020202020202020202020202020202020 //  net index:    34, net name:     n100                 
6e31303120202020202020202020202020202020 //  net index:    35, net name:     n101                 
6e31303220202020202020202020202020202020 //  net index:    36, net name:     n102                 
6e31303320202020202020202020202020202020 //  net index:    37, net name:     n103                 
6e31303420202020202020202020202020202020 //  net index:    38, net name:     n104                 
6e31303520202020202020202020202020202020 //  net index:    39, net name:     n105                 
6e31303620202020202020202020202020202020 //  net index:    40, net name:     n106                 
6e31303720202020202020202020202020202020 //  net index:    41, net name:     n107                 
6e31303820202020202020202020202020202020 //  net index:    42, net name:     n108                 
6e31303920202020202020202020202020202020 //  net index:    43, net name:     n109                 
6e31312020202020202020202020202020202020 //  net index:    44, net name:     n11                  
6e31313020202020202020202020202020202020 //  net index:    45, net name:     n110                 
6e31313120202020202020202020202020202020 //  net index:    46, net name:     n111                 
6e31313220202020202020202020202020202020 //  net index:    47, net name:     n112                 
6e31313320202020202020202020202020202020 //  net index:    48, net name:     n113                 
6e31313420202020202020202020202020202020 //  net index:    49, net name:     n114                 
6e31313520202020202020202020202020202020 //  net index:    50, net name:     n115                 
6e31313620202020202020202020202020202020 //  net index:    51, net name:     n116                 
6e31313720202020202020202020202020202020 //  net index:    52, net name:     n117                 
6e31313820202020202020202020202020202020 //  net index:    53, net name:     n118                 
6e31313920202020202020202020202020202020 //  net index:    54, net name:     n119                 
6e31322020202020202020202020202020202020 //  net index:    55, net name:     n12                  
6e31323020202020202020202020202020202020 //  net index:    56, net name:     n120                 
6e31323120202020202020202020202020202020 //  net index:    57, net name:     n121                 
6e31323220202020202020202020202020202020 //  net index:    58, net name:     n122                 
6e31323320202020202020202020202020202020 //  net index:    59, net name:     n123                 
6e31323420202020202020202020202020202020 //  net index:    60, net name:     n124                 
6e31323520202020202020202020202020202020 //  net index:    61, net name:     n125                 
6e31323620202020202020202020202020202020 //  net index:    62, net name:     n126                 
6e31323720202020202020202020202020202020 //  net index:    63, net name:     n127                 
6e31323820202020202020202020202020202020 //  net index:    64, net name:     n128                 
6e31323920202020202020202020202020202020 //  net index:    65, net name:     n129                 
6e31332020202020202020202020202020202020 //  net index:    66, net name:     n13                  
6e31333020202020202020202020202020202020 //  net index:    67, net name:     n130                 
6e31333120202020202020202020202020202020 //  net index:    68, net name:     n131                 
6e31333220202020202020202020202020202020 //  net index:    69, net name:     n132                 
6e31333320202020202020202020202020202020 //  net index:    70, net name:     n133                 
6e31333420202020202020202020202020202020 //  net index:    71, net name:     n134                 
6e31333520202020202020202020202020202020 //  net index:    72, net name:     n135                 
6e31333620202020202020202020202020202020 //  net index:    73, net name:     n136                 
6e31333720202020202020202020202020202020 //  net index:    74, net name:     n137                 
6e31333820202020202020202020202020202020 //  net index:    75, net name:     n138                 
6e31333920202020202020202020202020202020 //  net index:    76, net name:     n139                 
6e31342020202020202020202020202020202020 //  net index:    77, net name:     n14                  
6e31343020202020202020202020202020202020 //  net index:    78, net name:     n140                 
6e31343120202020202020202020202020202020 //  net index:    79, net name:     n141                 
6e31343220202020202020202020202020202020 //  net index:    80, net name:     n142                 
6e31343320202020202020202020202020202020 //  net index:    81, net name:     n143                 
6e31343420202020202020202020202020202020 //  net index:    82, net name:     n144                 
6e31343520202020202020202020202020202020 //  net index:    83, net name:     n145                 
6e31343620202020202020202020202020202020 //  net index:    84, net name:     n146                 
6e31343720202020202020202020202020202020 //  net index:    85, net name:     n147                 
6e31343820202020202020202020202020202020 //  net index:    86, net name:     n148                 
6e31343920202020202020202020202020202020 //  net index:    87, net name:     n149                 
6e31352020202020202020202020202020202020 //  net index:    88, net name:     n15                  
6e31353020202020202020202020202020202020 //  net index:    89, net name:     n150                 
6e31353120202020202020202020202020202020 //  net index:    90, net name:     n151                 
6e31353220202020202020202020202020202020 //  net index:    91, net name:     n152                 
6e31353320202020202020202020202020202020 //  net index:    92, net name:     n153                 
6e31353420202020202020202020202020202020 //  net index:    93, net name:     n154                 
6e31353520202020202020202020202020202020 //  net index:    94, net name:     n155                 
6e31353620202020202020202020202020202020 //  net index:    95, net name:     n156                 
6e31353720202020202020202020202020202020 //  net index:    96, net name:     n157                 
6e31353820202020202020202020202020202020 //  net index:    97, net name:     n158                 
6e31353920202020202020202020202020202020 //  net index:    98, net name:     n159                 
6e31362020202020202020202020202020202020 //  net index:    99, net name:     n16                  
6e31363020202020202020202020202020202020 //  net index:   100, net name:     n160                 
6e31363120202020202020202020202020202020 //  net index:   101, net name:     n161                 
6e31363220202020202020202020202020202020 //  net index:   102, net name:     n162                 
6e31363320202020202020202020202020202020 //  net index:   103, net name:     n163                 
6e31363420202020202020202020202020202020 //  net index:   104, net name:     n164                 
6e31372020202020202020202020202020202020 //  net index:   105, net name:     n17                  
6e31382020202020202020202020202020202020 //  net index:   106, net name:     n18                  
6e31392020202020202020202020202020202020 //  net index:   107, net name:     n19                  
6e32202020202020202020202020202020202020 //  net index:   108, net name:     n2                   
6e32302020202020202020202020202020202020 //  net index:   109, net name:     n20                  
6e32312020202020202020202020202020202020 //  net index:   110, net name:     n21                  
6e32322020202020202020202020202020202020 //  net index:   111, net name:     n22                  
6e32332020202020202020202020202020202020 //  net index:   112, net name:     n23                  
6e32342020202020202020202020202020202020 //  net index:   113, net name:     n24                  
6e32352020202020202020202020202020202020 //  net index:   114, net name:     n25                  
6e32362020202020202020202020202020202020 //  net index:   115, net name:     n26                  
6e32372020202020202020202020202020202020 //  net index:   116, net name:     n27                  
6e32382020202020202020202020202020202020 //  net index:   117, net name:     n28                  
6e32392020202020202020202020202020202020 //  net index:   118, net name:     n29                  
6e33202020202020202020202020202020202020 //  net index:   119, net name:     n3                   
6e33302020202020202020202020202020202020 //  net index:   120, net name:     n30                  
6e33312020202020202020202020202020202020 //  net index:   121, net name:     n31                  
6e33322020202020202020202020202020202020 //  net index:   122, net name:     n32                  
6e33332020202020202020202020202020202020 //  net index:   123, net name:     n33                  
6e33342020202020202020202020202020202020 //  net index:   124, net name:     n34                  
6e33352020202020202020202020202020202020 //  net index:   125, net name:     n35                  
6e33362020202020202020202020202020202020 //  net index:   126, net name:     n36                  
6e33372020202020202020202020202020202020 //  net index:   127, net name:     n37                  
6e33382020202020202020202020202020202020 //  net index:   128, net name:     n38                  
6e33392020202020202020202020202020202020 //  net index:   129, net name:     n39                  
6e34202020202020202020202020202020202020 //  net index:   130, net name:     n4                   
6e34302020202020202020202020202020202020 //  net index:   131, net name:     n40                  
6e34312020202020202020202020202020202020 //  net index:   132, net name:     n41                  
6e34322020202020202020202020202020202020 //  net index:   133, net name:     n42                  
6e34332020202020202020202020202020202020 //  net index:   134, net name:     n43                  
6e34342020202020202020202020202020202020 //  net index:   135, net name:     n44                  
6e34352020202020202020202020202020202020 //  net index:   136, net name:     n45                  
6e34362020202020202020202020202020202020 //  net index:   137, net name:     n46                  
6e34372020202020202020202020202020202020 //  net index:   138, net name:     n47                  
6e34382020202020202020202020202020202020 //  net index:   139, net name:     n48                  
6e34392020202020202020202020202020202020 //  net index:   140, net name:     n49                  
6e35202020202020202020202020202020202020 //  net index:   141, net name:     n5                   
6e35302020202020202020202020202020202020 //  net index:   142, net name:     n50                  
6e35312020202020202020202020202020202020 //  net index:   143, net name:     n51                  
6e35322020202020202020202020202020202020 //  net index:   144, net name:     n52                  
6e35332020202020202020202020202020202020 //  net index:   145, net name:     n53                  
6e35342020202020202020202020202020202020 //  net index:   146, net name:     n54                  
6e35352020202020202020202020202020202020 //  net index:   147, net name:     n55                  
6e35362020202020202020202020202020202020 //  net index:   148, net name:     n56                  
6e35372020202020202020202020202020202020 //  net index:   149, net name:     n57                  
6e35382020202020202020202020202020202020 //  net index:   150, net name:     n58                  
6e35392020202020202020202020202020202020 //  net index:   151, net name:     n59                  
6e36202020202020202020202020202020202020 //  net index:   152, net name:     n6                   
6e36302020202020202020202020202020202020 //  net index:   153, net name:     n60                  
6e36312020202020202020202020202020202020 //  net index:   154, net name:     n61                  
6e36322020202020202020202020202020202020 //  net index:   155, net name:     n62                  
6e36332020202020202020202020202020202020 //  net index:   156, net name:     n63                  
6e36342020202020202020202020202020202020 //  net index:   157, net name:     n64                  
6e36352020202020202020202020202020202020 //  net index:   158, net name:     n65                  
6e36362020202020202020202020202020202020 //  net index:   159, net name:     n66                  
6e36372020202020202020202020202020202020 //  net index:   160, net name:     n67                  
6e36382020202020202020202020202020202020 //  net index:   161, net name:     n68                  
6e36392020202020202020202020202020202020 //  net index:   162, net name:     n69                  
6e37202020202020202020202020202020202020 //  net index:   163, net name:     n7                   
6e37302020202020202020202020202020202020 //  net index:   164, net name:     n70                  
6e37312020202020202020202020202020202020 //  net index:   165, net name:     n71                  
6e37322020202020202020202020202020202020 //  net index:   166, net name:     n72                  
6e37332020202020202020202020202020202020 //  net index:   167, net name:     n73                  
6e37342020202020202020202020202020202020 //  net index:   168, net name:     n74                  
6e37352020202020202020202020202020202020 //  net index:   169, net name:     n75                  
6e37362020202020202020202020202020202020 //  net index:   170, net name:     n76                  
6e37372020202020202020202020202020202020 //  net index:   171, net name:     n77                  
6e37382020202020202020202020202020202020 //  net index:   172, net name:     n78                  
6e37392020202020202020202020202020202020 //  net index:   173, net name:     n79                  
6e38202020202020202020202020202020202020 //  net index:   174, net name:     n8                   
6e38302020202020202020202020202020202020 //  net index:   175, net name:     n80                  
6e38312020202020202020202020202020202020 //  net index:   176, net name:     n81                  
6e38322020202020202020202020202020202020 //  net index:   177, net name:     n82                  
6e38332020202020202020202020202020202020 //  net index:   178, net name:     n83                  
6e38342020202020202020202020202020202020 //  net index:   179, net name:     n84                  
6e38352020202020202020202020202020202020 //  net index:   180, net name:     n85                  
6e38362020202020202020202020202020202020 //  net index:   181, net name:     n86                  
6e38372020202020202020202020202020202020 //  net index:   182, net name:     n87                  
6e38382020202020202020202020202020202020 //  net index:   183, net name:     n88                  
6e38392020202020202020202020202020202020 //  net index:   184, net name:     n89                  
6e39202020202020202020202020202020202020 //  net index:   185, net name:     n9                   
6e39302020202020202020202020202020202020 //  net index:   186, net name:     n90                  
6e39312020202020202020202020202020202020 //  net index:   187, net name:     n91                  
6e39322020202020202020202020202020202020 //  net index:   188, net name:     n92                  
6e39332020202020202020202020202020202020 //  net index:   189, net name:     n93                  
6e39342020202020202020202020202020202020 //  net index:   190, net name:     n94                  
6e39352020202020202020202020202020202020 //  net index:   191, net name:     n95                  
6e39362020202020202020202020202020202020 //  net index:   192, net name:     n96                  
6e39372020202020202020202020202020202020 //  net index:   193, net name:     n97                  
6e39382020202020202020202020202020202020 //  net index:   194, net name:     n98                  
6e39392020202020202020202020202020202020 //  net index:   195, net name:     n99                  
6f5b305d20202020202020202020202020202020 //  net index:   196, net name:     o[0]                 output
6f5b31305d202020202020202020202020202020 //  net index:   197, net name:     o[10]                output
6f5b31315d202020202020202020202020202020 //  net index:   198, net name:     o[11]                output
6f5b31325d202020202020202020202020202020 //  net index:   199, net name:     o[12]                output
6f5b31335d202020202020202020202020202020 //  net index:   200, net name:     o[13]                output
6f5b31345d202020202020202020202020202020 //  net index:   201, net name:     o[14]                output
6f5b31355d202020202020202020202020202020 //  net index:   202, net name:     o[15]                output
6f5b315d20202020202020202020202020202020 //  net index:   203, net name:     o[1]                 output
6f5b325d20202020202020202020202020202020 //  net index:   204, net name:     o[2]                 output
6f5b335d20202020202020202020202020202020 //  net index:   205, net name:     o[3]                 output
6f5b345d20202020202020202020202020202020 //  net index:   206, net name:     o[4]                 output
6f5b355d20202020202020202020202020202020 //  net index:   207, net name:     o[5]                 output
6f5b365d20202020202020202020202020202020 //  net index:   208, net name:     o[6]                 output
6f5b375d20202020202020202020202020202020 //  net index:   209, net name:     o[7]                 output
6f5b385d20202020202020202020202020202020 //  net index:   210, net name:     o[8]                 output
6f5b395d20202020202020202020202020202020 //  net index:   211, net name:     o[9]                 output
