// DATA derived from module add1 !!!!!!!!!!!!!!!!
// code used to capture all changes in ref_dut and
// generates screen prints with time, value and net name
always @( ref_dut.a[0] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name a[0]",delta_time,ref_dut.a[0]); end
always @( ref_dut.a[10] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name a[10]",delta_time,ref_dut.a[10]); end
always @( ref_dut.a[11] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name a[11]",delta_time,ref_dut.a[11]); end
always @( ref_dut.a[12] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name a[12]",delta_time,ref_dut.a[12]); end
always @( ref_dut.a[13] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name a[13]",delta_time,ref_dut.a[13]); end
always @( ref_dut.a[14] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name a[14]",delta_time,ref_dut.a[14]); end
always @( ref_dut.a[15] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name a[15]",delta_time,ref_dut.a[15]); end
always @( ref_dut.a[1] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name a[1]",delta_time,ref_dut.a[1]); end
always @( ref_dut.a[2] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name a[2]",delta_time,ref_dut.a[2]); end
always @( ref_dut.a[3] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name a[3]",delta_time,ref_dut.a[3]); end
always @( ref_dut.a[4] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name a[4]",delta_time,ref_dut.a[4]); end
always @( ref_dut.a[5] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name a[5]",delta_time,ref_dut.a[5]); end
always @( ref_dut.a[6] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name a[6]",delta_time,ref_dut.a[6]); end
always @( ref_dut.a[7] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name a[7]",delta_time,ref_dut.a[7]); end
always @( ref_dut.a[8] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name a[8]",delta_time,ref_dut.a[8]); end
always @( ref_dut.a[9] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name a[9]",delta_time,ref_dut.a[9]); end
always @( ref_dut.b[0] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name b[0]",delta_time,ref_dut.b[0]); end
always @( ref_dut.b[10] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name b[10]",delta_time,ref_dut.b[10]); end
always @( ref_dut.b[11] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name b[11]",delta_time,ref_dut.b[11]); end
always @( ref_dut.b[12] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name b[12]",delta_time,ref_dut.b[12]); end
always @( ref_dut.b[13] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name b[13]",delta_time,ref_dut.b[13]); end
always @( ref_dut.b[14] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name b[14]",delta_time,ref_dut.b[14]); end
always @( ref_dut.b[15] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name b[15]",delta_time,ref_dut.b[15]); end
always @( ref_dut.b[1] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name b[1]",delta_time,ref_dut.b[1]); end
always @( ref_dut.b[2] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name b[2]",delta_time,ref_dut.b[2]); end
always @( ref_dut.b[3] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name b[3]",delta_time,ref_dut.b[3]); end
always @( ref_dut.b[4] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name b[4]",delta_time,ref_dut.b[4]); end
always @( ref_dut.b[5] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name b[5]",delta_time,ref_dut.b[5]); end
always @( ref_dut.b[6] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name b[6]",delta_time,ref_dut.b[6]); end
always @( ref_dut.b[7] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name b[7]",delta_time,ref_dut.b[7]); end
always @( ref_dut.b[8] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name b[8]",delta_time,ref_dut.b[8]); end
always @( ref_dut.b[9] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name b[9]",delta_time,ref_dut.b[9]); end
always @( ref_dut.n1 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n1",delta_time,ref_dut.n1); end
always @( ref_dut.n10 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n10",delta_time,ref_dut.n10); end
always @( ref_dut.n100 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n100",delta_time,ref_dut.n100); end
always @( ref_dut.n101 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n101",delta_time,ref_dut.n101); end
always @( ref_dut.n102 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n102",delta_time,ref_dut.n102); end
always @( ref_dut.n103 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n103",delta_time,ref_dut.n103); end
always @( ref_dut.n104 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n104",delta_time,ref_dut.n104); end
always @( ref_dut.n105 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n105",delta_time,ref_dut.n105); end
always @( ref_dut.n106 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n106",delta_time,ref_dut.n106); end
always @( ref_dut.n107 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n107",delta_time,ref_dut.n107); end
always @( ref_dut.n108 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n108",delta_time,ref_dut.n108); end
always @( ref_dut.n109 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n109",delta_time,ref_dut.n109); end
always @( ref_dut.n11 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n11",delta_time,ref_dut.n11); end
always @( ref_dut.n110 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n110",delta_time,ref_dut.n110); end
always @( ref_dut.n111 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n111",delta_time,ref_dut.n111); end
always @( ref_dut.n112 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n112",delta_time,ref_dut.n112); end
always @( ref_dut.n113 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n113",delta_time,ref_dut.n113); end
always @( ref_dut.n114 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n114",delta_time,ref_dut.n114); end
always @( ref_dut.n115 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n115",delta_time,ref_dut.n115); end
always @( ref_dut.n116 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n116",delta_time,ref_dut.n116); end
always @( ref_dut.n117 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n117",delta_time,ref_dut.n117); end
always @( ref_dut.n118 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n118",delta_time,ref_dut.n118); end
always @( ref_dut.n119 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n119",delta_time,ref_dut.n119); end
always @( ref_dut.n12 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n12",delta_time,ref_dut.n12); end
always @( ref_dut.n120 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n120",delta_time,ref_dut.n120); end
always @( ref_dut.n121 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n121",delta_time,ref_dut.n121); end
always @( ref_dut.n122 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n122",delta_time,ref_dut.n122); end
always @( ref_dut.n123 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n123",delta_time,ref_dut.n123); end
always @( ref_dut.n124 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n124",delta_time,ref_dut.n124); end
always @( ref_dut.n125 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n125",delta_time,ref_dut.n125); end
always @( ref_dut.n126 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n126",delta_time,ref_dut.n126); end
always @( ref_dut.n127 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n127",delta_time,ref_dut.n127); end
always @( ref_dut.n128 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n128",delta_time,ref_dut.n128); end
always @( ref_dut.n129 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n129",delta_time,ref_dut.n129); end
always @( ref_dut.n13 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n13",delta_time,ref_dut.n13); end
always @( ref_dut.n130 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n130",delta_time,ref_dut.n130); end
always @( ref_dut.n131 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n131",delta_time,ref_dut.n131); end
always @( ref_dut.n132 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n132",delta_time,ref_dut.n132); end
always @( ref_dut.n133 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n133",delta_time,ref_dut.n133); end
always @( ref_dut.n134 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n134",delta_time,ref_dut.n134); end
always @( ref_dut.n135 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n135",delta_time,ref_dut.n135); end
always @( ref_dut.n136 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n136",delta_time,ref_dut.n136); end
always @( ref_dut.n137 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n137",delta_time,ref_dut.n137); end
always @( ref_dut.n138 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n138",delta_time,ref_dut.n138); end
always @( ref_dut.n139 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n139",delta_time,ref_dut.n139); end
always @( ref_dut.n14 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n14",delta_time,ref_dut.n14); end
always @( ref_dut.n140 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n140",delta_time,ref_dut.n140); end
always @( ref_dut.n141 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n141",delta_time,ref_dut.n141); end
always @( ref_dut.n142 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n142",delta_time,ref_dut.n142); end
always @( ref_dut.n143 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n143",delta_time,ref_dut.n143); end
always @( ref_dut.n144 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n144",delta_time,ref_dut.n144); end
always @( ref_dut.n145 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n145",delta_time,ref_dut.n145); end
always @( ref_dut.n146 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n146",delta_time,ref_dut.n146); end
always @( ref_dut.n147 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n147",delta_time,ref_dut.n147); end
always @( ref_dut.n148 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n148",delta_time,ref_dut.n148); end
always @( ref_dut.n149 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n149",delta_time,ref_dut.n149); end
always @( ref_dut.n15 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n15",delta_time,ref_dut.n15); end
always @( ref_dut.n150 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n150",delta_time,ref_dut.n150); end
always @( ref_dut.n151 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n151",delta_time,ref_dut.n151); end
always @( ref_dut.n152 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n152",delta_time,ref_dut.n152); end
always @( ref_dut.n153 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n153",delta_time,ref_dut.n153); end
always @( ref_dut.n154 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n154",delta_time,ref_dut.n154); end
always @( ref_dut.n155 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n155",delta_time,ref_dut.n155); end
always @( ref_dut.n156 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n156",delta_time,ref_dut.n156); end
always @( ref_dut.n157 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n157",delta_time,ref_dut.n157); end
always @( ref_dut.n158 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n158",delta_time,ref_dut.n158); end
always @( ref_dut.n159 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n159",delta_time,ref_dut.n159); end
always @( ref_dut.n16 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n16",delta_time,ref_dut.n16); end
always @( ref_dut.n160 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n160",delta_time,ref_dut.n160); end
always @( ref_dut.n161 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n161",delta_time,ref_dut.n161); end
always @( ref_dut.n162 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n162",delta_time,ref_dut.n162); end
always @( ref_dut.n163 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n163",delta_time,ref_dut.n163); end
always @( ref_dut.n164 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n164",delta_time,ref_dut.n164); end
always @( ref_dut.n17 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n17",delta_time,ref_dut.n17); end
always @( ref_dut.n18 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n18",delta_time,ref_dut.n18); end
always @( ref_dut.n19 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n19",delta_time,ref_dut.n19); end
always @( ref_dut.n2 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n2",delta_time,ref_dut.n2); end
always @( ref_dut.n20 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n20",delta_time,ref_dut.n20); end
always @( ref_dut.n21 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n21",delta_time,ref_dut.n21); end
always @( ref_dut.n22 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n22",delta_time,ref_dut.n22); end
always @( ref_dut.n23 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n23",delta_time,ref_dut.n23); end
always @( ref_dut.n24 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n24",delta_time,ref_dut.n24); end
always @( ref_dut.n25 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n25",delta_time,ref_dut.n25); end
always @( ref_dut.n26 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n26",delta_time,ref_dut.n26); end
always @( ref_dut.n27 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n27",delta_time,ref_dut.n27); end
always @( ref_dut.n28 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n28",delta_time,ref_dut.n28); end
always @( ref_dut.n29 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n29",delta_time,ref_dut.n29); end
always @( ref_dut.n3 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n3",delta_time,ref_dut.n3); end
always @( ref_dut.n30 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n30",delta_time,ref_dut.n30); end
always @( ref_dut.n31 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n31",delta_time,ref_dut.n31); end
always @( ref_dut.n32 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n32",delta_time,ref_dut.n32); end
always @( ref_dut.n33 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n33",delta_time,ref_dut.n33); end
always @( ref_dut.n34 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n34",delta_time,ref_dut.n34); end
always @( ref_dut.n35 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n35",delta_time,ref_dut.n35); end
always @( ref_dut.n36 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n36",delta_time,ref_dut.n36); end
always @( ref_dut.n37 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n37",delta_time,ref_dut.n37); end
always @( ref_dut.n38 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n38",delta_time,ref_dut.n38); end
always @( ref_dut.n39 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n39",delta_time,ref_dut.n39); end
always @( ref_dut.n4 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n4",delta_time,ref_dut.n4); end
always @( ref_dut.n40 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n40",delta_time,ref_dut.n40); end
always @( ref_dut.n41 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n41",delta_time,ref_dut.n41); end
always @( ref_dut.n42 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n42",delta_time,ref_dut.n42); end
always @( ref_dut.n43 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n43",delta_time,ref_dut.n43); end
always @( ref_dut.n44 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n44",delta_time,ref_dut.n44); end
always @( ref_dut.n45 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n45",delta_time,ref_dut.n45); end
always @( ref_dut.n46 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n46",delta_time,ref_dut.n46); end
always @( ref_dut.n47 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n47",delta_time,ref_dut.n47); end
always @( ref_dut.n48 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n48",delta_time,ref_dut.n48); end
always @( ref_dut.n49 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n49",delta_time,ref_dut.n49); end
always @( ref_dut.n5 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n5",delta_time,ref_dut.n5); end
always @( ref_dut.n50 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n50",delta_time,ref_dut.n50); end
always @( ref_dut.n51 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n51",delta_time,ref_dut.n51); end
always @( ref_dut.n52 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n52",delta_time,ref_dut.n52); end
always @( ref_dut.n53 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n53",delta_time,ref_dut.n53); end
always @( ref_dut.n54 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n54",delta_time,ref_dut.n54); end
always @( ref_dut.n55 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n55",delta_time,ref_dut.n55); end
always @( ref_dut.n56 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n56",delta_time,ref_dut.n56); end
always @( ref_dut.n57 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n57",delta_time,ref_dut.n57); end
always @( ref_dut.n58 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n58",delta_time,ref_dut.n58); end
always @( ref_dut.n59 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n59",delta_time,ref_dut.n59); end
always @( ref_dut.n6 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n6",delta_time,ref_dut.n6); end
always @( ref_dut.n60 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n60",delta_time,ref_dut.n60); end
always @( ref_dut.n61 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n61",delta_time,ref_dut.n61); end
always @( ref_dut.n62 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n62",delta_time,ref_dut.n62); end
always @( ref_dut.n63 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n63",delta_time,ref_dut.n63); end
always @( ref_dut.n64 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n64",delta_time,ref_dut.n64); end
always @( ref_dut.n65 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n65",delta_time,ref_dut.n65); end
always @( ref_dut.n66 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n66",delta_time,ref_dut.n66); end
always @( ref_dut.n67 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n67",delta_time,ref_dut.n67); end
always @( ref_dut.n68 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n68",delta_time,ref_dut.n68); end
always @( ref_dut.n69 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n69",delta_time,ref_dut.n69); end
always @( ref_dut.n7 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n7",delta_time,ref_dut.n7); end
always @( ref_dut.n70 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n70",delta_time,ref_dut.n70); end
always @( ref_dut.n71 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n71",delta_time,ref_dut.n71); end
always @( ref_dut.n72 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n72",delta_time,ref_dut.n72); end
always @( ref_dut.n73 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n73",delta_time,ref_dut.n73); end
always @( ref_dut.n74 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n74",delta_time,ref_dut.n74); end
always @( ref_dut.n75 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n75",delta_time,ref_dut.n75); end
always @( ref_dut.n76 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n76",delta_time,ref_dut.n76); end
always @( ref_dut.n77 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n77",delta_time,ref_dut.n77); end
always @( ref_dut.n78 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n78",delta_time,ref_dut.n78); end
always @( ref_dut.n79 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n79",delta_time,ref_dut.n79); end
always @( ref_dut.n8 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n8",delta_time,ref_dut.n8); end
always @( ref_dut.n80 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n80",delta_time,ref_dut.n80); end
always @( ref_dut.n81 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n81",delta_time,ref_dut.n81); end
always @( ref_dut.n82 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n82",delta_time,ref_dut.n82); end
always @( ref_dut.n83 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n83",delta_time,ref_dut.n83); end
always @( ref_dut.n84 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n84",delta_time,ref_dut.n84); end
always @( ref_dut.n85 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n85",delta_time,ref_dut.n85); end
always @( ref_dut.n86 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n86",delta_time,ref_dut.n86); end
always @( ref_dut.n87 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n87",delta_time,ref_dut.n87); end
always @( ref_dut.n88 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n88",delta_time,ref_dut.n88); end
always @( ref_dut.n89 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n89",delta_time,ref_dut.n89); end
always @( ref_dut.n9 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n9",delta_time,ref_dut.n9); end
always @( ref_dut.n90 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n90",delta_time,ref_dut.n90); end
always @( ref_dut.n91 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n91",delta_time,ref_dut.n91); end
always @( ref_dut.n92 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n92",delta_time,ref_dut.n92); end
always @( ref_dut.n93 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n93",delta_time,ref_dut.n93); end
always @( ref_dut.n94 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n94",delta_time,ref_dut.n94); end
always @( ref_dut.n95 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n95",delta_time,ref_dut.n95); end
always @( ref_dut.n96 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n96",delta_time,ref_dut.n96); end
always @( ref_dut.n97 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n97",delta_time,ref_dut.n97); end
always @( ref_dut.n98 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n98",delta_time,ref_dut.n98); end
always @( ref_dut.n99 )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name n99",delta_time,ref_dut.n99); end
always @( ref_dut.o[0] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name o[0]",delta_time,ref_dut.o[0]); end
always @( ref_dut.o[10] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name o[10]",delta_time,ref_dut.o[10]); end
always @( ref_dut.o[11] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name o[11]",delta_time,ref_dut.o[11]); end
always @( ref_dut.o[12] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name o[12]",delta_time,ref_dut.o[12]); end
always @( ref_dut.o[13] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name o[13]",delta_time,ref_dut.o[13]); end
always @( ref_dut.o[14] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name o[14]",delta_time,ref_dut.o[14]); end
always @( ref_dut.o[15] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name o[15]",delta_time,ref_dut.o[15]); end
always @( ref_dut.o[1] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name o[1]",delta_time,ref_dut.o[1]); end
always @( ref_dut.o[2] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name o[2]",delta_time,ref_dut.o[2]); end
always @( ref_dut.o[3] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name o[3]",delta_time,ref_dut.o[3]); end
always @( ref_dut.o[4] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name o[4]",delta_time,ref_dut.o[4]); end
always @( ref_dut.o[5] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name o[5]",delta_time,ref_dut.o[5]); end
always @( ref_dut.o[6] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name o[6]",delta_time,ref_dut.o[6]); end
always @( ref_dut.o[7] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name o[7]",delta_time,ref_dut.o[7]); end
always @( ref_dut.o[8] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name o[8]",delta_time,ref_dut.o[8]); end
always @( ref_dut.o[9] )
	begin delta_time=($time-start_time); $display("===  ref_vcd      time %d ps, value %b, net name o[9]",delta_time,ref_dut.o[9]); end
