// DATA derived from module simple0 !!!!!!!!!!!!!!!!
// table used by testbench to translate out_records
// from turbosim to screen prints with time, value and net name
6120202020202020202020202020202020202020 //  net index:     0, net name:     a                    input
6220202020202020202020202020202020202020 //  net index:     1, net name:     b                    input
6320202020202020202020202020202020202020 //  net index:     2, net name:     c                    input
6420202020202020202020202020202020202020 //  net index:     3, net name:     d                    input
6520202020202020202020202020202020202020 //  net index:     4, net name:     e                    
6620202020202020202020202020202020202020 //  net index:     5, net name:     f                    
6720202020202020202020202020202020202020 //  net index:     6, net name:     g                    
6a31202020202020202020202020202020202020 //  net index:     7, net name:     j1                   
6a32202020202020202020202020202020202020 //  net index:     8, net name:     j2                   
6a33202020202020202020202020202020202020 //  net index:     9, net name:     j3                   
6e31202020202020202020202020202020202020 //  net index:    10, net name:     n1                   
6f31202020202020202020202020202020202020 //  net index:    11, net name:     o1                   output
6f32202020202020202020202020202020202020 //  net index:    12, net name:     o2                   output
