// DATA derived from module latch0 !!!!!!!!!!!!!!!!
// table used by testbench to translate out_records
// from turbosim to screen prints with time, value and net name
636c6b2020202020202020202020202020202020 //  net index:     0, net name:     clk                  input
6420202020202020202020202020202020202020 //  net index:     1, net name:     d                    input
6e31202020202020202020202020202020202020 //  net index:     2, net name:     n1                   
6e32202020202020202020202020202020202020 //  net index:     3, net name:     n2                   
6e33202020202020202020202020202020202020 //  net index:     4, net name:     n3                   
6e34202020202020202020202020202020202020 //  net index:     5, net name:     n4                   
6e35202020202020202020202020202020202020 //  net index:     6, net name:     n5                   
7120202020202020202020202020202020202020 //  net index:     7, net name:     q                    output
7162202020202020202020202020202020202020 //  net index:     8, net name:     qb                   output
